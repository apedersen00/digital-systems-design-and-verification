//-------------------------------------------------------------------------------------------------
//
//  File: cpu_pkg.sv
//  Description: Parameters and enums for CPU.
//
//  Author:
//      - A. Pedersen
//      - J. Sadiq
//      - J. Yang
//
//-------------------------------------------------------------------------------------------------

package core_pkg;

  `define 7'b0110011 R_INST
  `define 7'b

endpackage