//-------------------------------------------------------------------------------------------------
//
//  File: bin2gray.sv
//  Description: 4-bit binary to gray encoder.
//
//  Author:
//      - A. Pedersen
//
//-------------------------------------------------------------------------------------------------

//  bin2gray dut (
//    .binary(),
//    .gray()
//  );

module bin2gray (
    input   logic [3:0] binary,
    output  logic [3:0] gray
  );

  logic [15:0] gray_1_table = '{
    1'b0, // 1111
    0'b1, // 1110
    1'b1, // 1101
    0'b0, // 1100
    1'b0, // 1011
    0'b1, // 1010
    1'b1, // 1001
    0'b0, // 1000
    1'b0, // 0111
    0'b1, // 0110
    1'b1, // 0101
    0'b0, // 0100
    1'b0, // 0011
    0'b1, // 0010
    1'b1, // 0001
    0'b0  // 0000
  };

  logic [15:0] gray_2_table = '{
    1'b0, // 1111
    0'b0, // 1110
    1'b1, // 1101
    0'b1, // 1100
    1'b1, // 1011
    0'b1, // 1010
    1'b0, // 1001
    0'b0, // 1000
    1'b0, // 0111
    0'b0, // 0110
    1'b1, // 0101
    0'b1, // 0100
    1'b1, // 0011
    0'b1, // 0010
    1'b0, // 0001
    0'b0  // 0000
  };

  logic [15:0] gray_4_table = '{
    1'b0, // 1111
    0'b0, // 1110
    1'b0, // 1101
    0'b0, // 1100
    1'b1, // 1011
    0'b1, // 1010
    1'b1, // 1001
    0'b1, // 1000
    1'b1, // 0111
    0'b1, // 0110
    1'b1, // 0101
    0'b1, // 0100
    1'b0, // 0011
    0'b0, // 0010
    1'b0, // 0001
    0'b0  // 0000
  };

  logic [15:0] gray_8_table = '{
    1'b1, // 1111
    0'b1, // 1110
    1'b1, // 1101
    0'b1, // 1100
    1'b1, // 1011
    0'b1, // 1010
    1'b1, // 1001
    0'b1, // 1000
    1'b0, // 0111
    0'b0, // 0110
    1'b0, // 0101
    0'b0, // 0100
    1'b0, // 0011
    0'b0, // 0010
    1'b0, // 0001
    0'b0  // 0000
  };

  mux #(
    .InputWidth(16)
  ) mux_gray_1 (
    .in(gray_1_table),
    .select(binary),
    .out(gray[0])
  );

  mux #(
    .InputWidth(16)
  ) mux_gray_2 (
    .in(gray_2_table),
    .select(binary),
    .out(gray[1])
  );

  mux #(
    .InputWidth(16)
  ) mux_gray_4 (
    .in(gray_4_table),
    .select(binary),
    .out(gray[2])
  );

  mux #(
    .InputWidth(16)
  ) mux_gray_8 (
    .in(gray_8_table),
    .select(binary),
    .out(gray[3])
  );

endmodule