//-------------------------------------------------------------------------------------------------
//
//  File: reciprocal.sv
//  Description:
//
//  Author:
//
//-------------------------------------------------------------------------------------------------

//  reciprocal reciprocal_0 (
//    .x_i(),
//    .y_o()
//  );

module reciprocal ( 
    input  logic [15:0] x_i, 
    output logic [8:0]  y_o
  );
    
  always_comb begin
    case (x_i)
      16'h0001: y_o = 9'h100;   // 1
      16'h0002: y_o = 9'h080;   // 1/2
      16'h0003: y_o = 9'h055;   // 1/3
      16'h0004: y_o = 9'h040;   // 1/4
      16'h0005: y_o = 9'h033;   // 1/5
      16'h0006: y_o = 9'h02A;   // 1/6
      16'h0007: y_o = 9'h024;   // 1/7
      16'h0008: y_o = 9'h020;   // 1/8
      16'h0009: y_o = 9'h01C;   // 1/9
      16'h000A: y_o = 9'h019;   // 1/10
      16'h000B: y_o = 9'h017;   // 1/11
      16'h000C: y_o = 9'h015;   // 1/12
      16'h000D: y_o = 9'h013;   // 1/13
      16'h000E: y_o = 9'h012;   // 1/14
      16'h000F: y_o = 9'h011;   // 1/15
      default:  y_o = 9'h000;   // out of range, return 0
    endcase
  end

endmodule